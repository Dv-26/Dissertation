
module HuffmanCoder #(
parameter CHROMA = 1
) (
input logic clk, rst_n,
input tempCode_t in,
);
  localparam CODE_W = CHROMA == 1 ? 9 : 11;
  struct {
    logic [CODE_W-1:0] code,
    logic [3:0] size
  } DCHuffman;
  AcHuffman_t ACHuffman;

  DCHuffmanMap #(CHROMA) DCHuffmanMap (
    clk,
    in.data.size, in.data.isDC & in.valid,
    DCHuffman.code, DCHuffman.size
  );

  ACHuffmanMap #(CHROMA) ACHuffmanMap (
    clk,
    in.data.run, in.data.size, ~in.data.isDC & in.valid,
    ACHuffman
  );

endmodule

module DCHuffmanMap#(
  parameter CHROMA = 1
) (
  clk,
  size, en,
  huffmanCode, huffmanSize
);
  localparam CODE_W = CHROMA == 1 ? 9 : 11;

  input logic clk;
  input logic [$bits(tempCodeData_t.size)-1:0] size;
  input logic en;
  output logic [CODE_W-1:0] huffmanCode; 
  output logic [3:0] huffmanSize;

  always_ff @(posedge clk) begin
    if(en)
      {huffmanSize, huffmanCode} <= 
  end
  logic [CODE_W+$bits(huffmanSize)-1:0] array [12];
  initial begin
    if(CHROMA=1) begin
      array[4'h0] = {4'h2, 9'b000000000};
      array[4'h1] = {4'h3, 9'b000000010};
      array[4'h2] = {4'h3, 9'b000000011};
      array[4'h3] = {4'h3, 9'b000000100};
      array[4'h4] = {4'h3, 9'b000000101};
      array[4'h5] = {4'h3, 9'b000000110};
      array[4'h6] = {4'h4, 9'b000001110};
      array[4'h7] = {4'h5, 9'b000011110};
      array[4'h8] = {4'h6, 9'b000111110};
      array[4'h9] = {4'h7, 9'b001111110};
      array[4'ha] = {4'h9, 9'b011111110};
      array[4'hb] = {4'h9, 9'b111111110};
    end else begin
      array[4'h0] = {4'h2, 11'b00000000000};
      array[4'h1] = {4'h2, 11'b00000000001};
      array[4'h2] = {4'h2, 11'b00000000010};
      array[4'h3] = {4'h3, 11'b00000000110};
      array[4'h4] = {4'h4, 11'b00000001110};
      array[4'h5] = {4'h5, 11'b00000011110};
      array[4'h6] = {4'h6, 11'b00000111110};
      array[4'h7] = {4'h7, 11'b00001111110};
      array[4'h8] = {4'h8, 11'b00011111110};
      array[4'h9] = {4'h9, 11'b00111111110};
      array[4'ha] = {4'ha, 11'b01111111110};
      array[4'hb] = {4'hb, 11'b11111111110};
    end
  end
  
endmodule


module ACHuffmanMap#(
  parameter CHROMA = 1
) (
  clk,
  run, size, en,
  huffman
);
  input logic clk;
  input logic [$bits(tempCodeData_t.run)-1:0] run;
  input logic [$bits(tempCodeData_t.size)-1:0] size;
  input logic en;
  output AcHuffman_t huffman;

  logic [$bits(chrominanceAcHuffman_t)-1:0] array [162];
  always_ff @(posedge clk)
    if(en) 
      {huffman.size, huffman.code} <= array[{run, size}];

  initial begin
    if(CHROMA == 1) begin
      array[{4'h0, 4'h0}] = {5'd4, 16'b0000000000001010};
      array[{4'h0, 4'h1}] = {5'd2, 16'b0000000000000000};
      array[{4'h0, 4'h2}] = {5'd2, 16'b0000000000000001};
      array[{4'h0, 4'h3}] = {5'd3, 16'b0000000000000100};
      array[{4'h0, 4'h4}] = {5'd4, 16'b0000000000001011};
      array[{4'h0, 4'h5}] = {5'd5, 16'b0000000000011010};
      array[{4'h0, 4'h6}] = {5'd7, 16'b0000000001111000};
      array[{4'h0, 4'h7}] = {5'd8, 16'b0000000011111000};
      array[{4'h0, 4'h8}] = {5'd10, 16'b0000001111110110};
      array[{4'h0, 4'h9}] = {5'd16, 16'b1111111110000010};
      array[{4'h0, 4'hA}] = {5'd16, 16'b1111111110000011};
      array[{4'h1, 4'h1}] = {5'd4, 16'b0000000000001100};
      array[{4'h1, 4'h2}] = {5'd5, 16'b0000000000011011};
      array[{4'h1, 4'h3}] = {5'd7, 16'b0000000001111001};
      array[{4'h1, 4'h4}] = {5'd9, 16'b0000000111110110};
      array[{4'h1, 4'h5}] = {5'd11, 16'b0000011111110110};
      array[{4'h1, 4'h6}] = {5'd16, 16'b1111111110000100};
      array[{4'h1, 4'h7}] = {5'd16, 16'b1111111110000101};
      array[{4'h1, 4'h8}] = {5'd16, 16'b1111111110000110};
      array[{4'h1, 4'h9}] = {5'd16, 16'b1111111110000111};
      array[{4'h1, 4'hA}] = {5'd16, 16'b1111111110001000};
      array[{4'h2, 4'h1}] = {5'd5, 16'b0000000000011100};
      array[{4'h2, 4'h2}] = {5'd8, 16'b0000000011111001};
      array[{4'h2, 4'h3}] = {5'd10, 16'b0000001111110111};
      array[{4'h2, 4'h4}] = {5'd12, 16'b0000111111110100};
      array[{4'h2, 4'h5}] = {5'd16, 16'b1111111110001001};
      array[{4'h2, 4'h6}] = {5'd16, 16'b1111111110001010};
      array[{4'h2, 4'h7}] = {5'd16, 16'b1111111110001011};
      array[{4'h2, 4'h8}] = {5'd16, 16'b1111111110001100};
      array[{4'h2, 4'h9}] = {5'd16, 16'b1111111110001101};
      array[{4'h2, 4'hA}] = {5'd16, 16'b1111111110001110};
      array[{4'h3, 4'h1}] = {5'd6, 16'b0000000000111010};
      array[{4'h3, 4'h2}] = {5'd9, 16'b0000000111110111};
      array[{4'h3, 4'h3}] = {5'd12, 16'b0000111111110101};
      array[{4'h3, 4'h4}] = {5'd16, 16'b1111111110001111};
      array[{4'h3, 4'h5}] = {5'd16, 16'b1111111110010000};
      array[{4'h3, 4'h6}] = {5'd16, 16'b1111111110010001};
      array[{4'h3, 4'h7}] = {5'd16, 16'b1111111110010010};
      array[{4'h3, 4'h8}] = {5'd16, 16'b1111111110010011};
      array[{4'h3, 4'h9}] = {5'd16, 16'b1111111110010100};
      array[{4'h3, 4'hA}] = {5'd16, 16'b1111111110010101};
      array[{4'h4, 4'h1}] = {5'd6, 16'b0000000000111011};
      array[{4'h4, 4'h2}] = {5'd10, 16'b0000001111111000};
      array[{4'h4, 4'h3}] = {5'd16, 16'b1111111110010110};
      array[{4'h4, 4'h4}] = {5'd16, 16'b1111111110010111};
      array[{4'h4, 4'h5}] = {5'd16, 16'b1111111110011000};
      array[{4'h4, 4'h6}] = {5'd16, 16'b1111111110011001};
      array[{4'h4, 4'h7}] = {5'd16, 16'b1111111110011010};
      array[{4'h4, 4'h8}] = {5'd16, 16'b1111111110011011};
      array[{4'h4, 4'h9}] = {5'd16, 16'b1111111110011100};
      array[{4'h4, 4'hA}] = {5'd16, 16'b1111111110011101};
      array[{4'h5, 4'h1}] = {5'd7, 16'b0000000001111010};
      array[{4'h5, 4'h2}] = {5'd11, 16'b0000011111110111};
      array[{4'h5, 4'h3}] = {5'd16, 16'b1111111110011110};
      array[{4'h5, 4'h4}] = {5'd16, 16'b1111111110011111};
      array[{4'h5, 4'h5}] = {5'd16, 16'b1111111110100000};
      array[{4'h5, 4'h6}] = {5'd16, 16'b1111111110100001};
      array[{4'h5, 4'h7}] = {5'd16, 16'b1111111110100010};
      array[{4'h5, 4'h8}] = {5'd16, 16'b1111111110100011};
      array[{4'h5, 4'h9}] = {5'd16, 16'b1111111110100100};
      array[{4'h5, 4'hA}] = {5'd16, 16'b1111111110100101};
      array[{4'h6, 4'h1}] = {5'd7, 16'b0000000001111011};
      array[{4'h6, 4'h2}] = {5'd12, 16'b0000111111110110};
      array[{4'h6, 4'h3}] = {5'd16, 16'b1111111110100110};
      array[{4'h6, 4'h4}] = {5'd16, 16'b1111111110100111};
      array[{4'h6, 4'h5}] = {5'd16, 16'b1111111110101000};
      array[{4'h6, 4'h6}] = {5'd16, 16'b1111111110101001};
      array[{4'h6, 4'h7}] = {5'd16, 16'b1111111110101010};
      array[{4'h6, 4'h8}] = {5'd16, 16'b1111111110101011};
      array[{4'h6, 4'h9}] = {5'd16, 16'b1111111110101100};
      array[{4'h6, 4'hA}] = {5'd16, 16'b1111111110101101};
      array[{4'h7, 4'h1}] = {5'd8, 16'b0000000011111010};
      array[{4'h7, 4'h2}] = {5'd12, 16'b0000111111110111};
      array[{4'h7, 4'h3}] = {5'd16, 16'b1111111110101110};
      array[{4'h7, 4'h4}] = {5'd16, 16'b1111111110101111};
      array[{4'h7, 4'h5}] = {5'd16, 16'b1111111110110000};
      array[{4'h7, 4'h6}] = {5'd16, 16'b1111111110110001};
      array[{4'h7, 4'h7}] = {5'd16, 16'b1111111110110010};
      array[{4'h7, 4'h8}] = {5'd16, 16'b1111111110110011};
      array[{4'h7, 4'h9}] = {5'd16, 16'b1111111110110100};
      array[{4'h7, 4'hA}] = {5'd16, 16'b1111111110110101};
      array[{4'h8, 4'h1}] = {5'd9, 16'b0000000111111000};
      array[{4'h8, 4'h2}] = {5'd15, 16'b0111111111000000};
      array[{4'h8, 4'h3}] = {5'd16, 16'b1111111110110110};
      array[{4'h8, 4'h4}] = {5'd16, 16'b1111111110110111};
      array[{4'h8, 4'h5}] = {5'd16, 16'b1111111110111000};
      array[{4'h8, 4'h6}] = {5'd16, 16'b1111111110111001};
      array[{4'h8, 4'h7}] = {5'd16, 16'b1111111110111010};
      array[{4'h8, 4'h8}] = {5'd16, 16'b1111111110111011};
      array[{4'h8, 4'h9}] = {5'd16, 16'b1111111110111100};
      array[{4'h8, 4'hA}] = {5'd16, 16'b1111111110111101};
      array[{4'h9, 4'h1}] = {5'd9, 16'b0000000111111001};
      array[{4'h9, 4'h2}] = {5'd16, 16'b1111111110111110};
      array[{4'h9, 4'h3}] = {5'd16, 16'b1111111110111111};
      array[{4'h9, 4'h4}] = {5'd16, 16'b1111111111000000};
      array[{4'h9, 4'h5}] = {5'd16, 16'b1111111111000001};
      array[{4'h9, 4'h6}] = {5'd16, 16'b1111111111000010};
      array[{4'h9, 4'h7}] = {5'd16, 16'b1111111111000011};
      array[{4'h9, 4'h8}] = {5'd16, 16'b1111111111000100};
      array[{4'h9, 4'h9}] = {5'd16, 16'b1111111111000101};
      array[{4'h9, 4'hA}] = {5'd16, 16'b1111111111000110};
      array[{4'hA, 4'h1}] = {5'd9, 16'b0000000111111010};
      array[{4'hA, 4'h2}] = {5'd16, 16'b1111111111000111};
      array[{4'hA, 4'h3}] = {5'd16, 16'b1111111111001000};
      array[{4'hA, 4'h4}] = {5'd16, 16'b1111111111001001};
      array[{4'hA, 4'h5}] = {5'd16, 16'b1111111111001010};
      array[{4'hA, 4'h6}] = {5'd16, 16'b1111111111001011};
      array[{4'hA, 4'h7}] = {5'd16, 16'b1111111111001100};
      array[{4'hA, 4'h8}] = {5'd16, 16'b1111111111001101};
      array[{4'hA, 4'h9}] = {5'd16, 16'b1111111111001110};
      array[{4'hA, 4'hA}] = {5'd16, 16'b1111111111001111};
      array[{4'hB, 4'h1}] = {5'd10, 16'b0000001111111001};
      array[{4'hB, 4'h2}] = {5'd16, 16'b1111111111010000};
      array[{4'hB, 4'h3}] = {5'd16, 16'b1111111111010001};
      array[{4'hB, 4'h4}] = {5'd16, 16'b1111111111010010};
      array[{4'hB, 4'h5}] = {5'd16, 16'b1111111111010011};
      array[{4'hB, 4'h6}] = {5'd16, 16'b1111111111010100};
      array[{4'hB, 4'h7}] = {5'd16, 16'b1111111111010101};
      array[{4'hB, 4'h8}] = {5'd16, 16'b1111111111010110};
      array[{4'hB, 4'h9}] = {5'd16, 16'b1111111111010111};
      array[{4'hB, 4'hA}] = {5'd16, 16'b1111111111011000};
      array[{4'hC, 4'h1}] = {5'd10, 16'b0000001111111010};
      array[{4'hC, 4'h2}] = {5'd16, 16'b1111111111011001};
      array[{4'hC, 4'h3}] = {5'd16, 16'b1111111111011010};
      array[{4'hC, 4'h4}] = {5'd16, 16'b1111111111011011};
      array[{4'hC, 4'h5}] = {5'd16, 16'b1111111111011100};
      array[{4'hC, 4'h6}] = {5'd16, 16'b1111111111011101};
      array[{4'hC, 4'h7}] = {5'd16, 16'b1111111111011110};
      array[{4'hC, 4'h8}] = {5'd16, 16'b1111111111011111};
      array[{4'hC, 4'h9}] = {5'd16, 16'b1111111111100000};
      array[{4'hC, 4'hA}] = {5'd16, 16'b1111111111100001};
      array[{4'hD, 4'h1}] = {5'd11, 16'b0000011111111000};
      array[{4'hD, 4'h2}] = {5'd16, 16'b1111111111100010};
      array[{4'hD, 4'h3}] = {5'd16, 16'b1111111111100011};
      array[{4'hD, 4'h4}] = {5'd16, 16'b1111111111100100};
      array[{4'hD, 4'h5}] = {5'd16, 16'b1111111111100101};
      array[{4'hD, 4'h6}] = {5'd16, 16'b1111111111100110};
      array[{4'hD, 4'h7}] = {5'd16, 16'b1111111111100111};
      array[{4'hD, 4'h8}] = {5'd16, 16'b1111111111101000};
      array[{4'hD, 4'h9}] = {5'd16, 16'b1111111111101001};
      array[{4'hD, 4'hA}] = {5'd16, 16'b1111111111101010};
      array[{4'hE, 4'h1}] = {5'd16, 16'b1111111111101011};
      array[{4'hE, 4'h2}] = {5'd16, 16'b1111111111101100};
      array[{4'hE, 4'h3}] = {5'd16, 16'b1111111111101101};
      array[{4'hE, 4'h4}] = {5'd16, 16'b1111111111101110};
      array[{4'hE, 4'h5}] = {5'd16, 16'b1111111111101111};
      array[{4'hE, 4'h6}] = {5'd16, 16'b1111111111110000};
      array[{4'hE, 4'h7}] = {5'd16, 16'b1111111111110001};
      array[{4'hE, 4'h8}] = {5'd16, 16'b1111111111110010};
      array[{4'hE, 4'h9}] = {5'd16, 16'b1111111111110011};
      array[{4'hE, 4'hA}] = {5'd16, 16'b1111111111110100};
      array[{4'hF, 4'h0}] = {5'd11, 16'b0000011111111001};
      array[{4'hF, 4'h1}] = {5'd16, 16'b1111111111110101};
      array[{4'hF, 4'h2}] = {5'd16, 16'b1111111111110110};
      array[{4'hF, 4'h3}] = {5'd16, 16'b1111111111110111};
      array[{4'hF, 4'h4}] = {5'd16, 16'b1111111111111000};
      array[{4'hF, 4'h5}] = {5'd16, 16'b1111111111111001};
      array[{4'hF, 4'h6}] = {5'd16, 16'b1111111111111010};
      array[{4'hF, 4'h7}] = {5'd16, 16'b1111111111111011};
      array[{4'hF, 4'h8}] = {5'd16, 16'b1111111111111100};
      array[{4'hF, 4'h9}] = {5'd16, 16'b1111111111111101};
      array[{4'hF, 4'hA}] = {5'd16, 16'b1111111111111110};
    end else begin
      array[{4'h0, 4'h0}] = {5'd2, 16'b0000000000000000};
      array[{4'h0, 4'h1}] = {5'd2, 16'b0000000000000001};
      array[{4'h0, 4'h2}] = {5'd3, 16'b0000000000000100};
      array[{4'h0, 4'h3}] = {5'd4, 16'b0000000000001010};
      array[{4'h0, 4'h4}] = {5'd5, 16'b0000000000011000};
      array[{4'h0, 4'h5}] = {5'd5, 16'b0000000000011001};
      array[{4'h0, 4'h6}] = {5'd6, 16'b0000000000111000};
      array[{4'h0, 4'h7}] = {5'd7, 16'b0000000001111000};
      array[{4'h0, 4'h8}] = {5'd9, 16'b0000000111110100};
      array[{4'h0, 4'h9}] = {5'd10, 16'b0000001111110110};
      array[{4'h0, 4'hA}] = {5'd12, 16'b0000111111110100};
      array[{4'h1, 4'h1}] = {5'd4, 16'b0000000000001011};
      array[{4'h1, 4'h2}] = {5'd6, 16'b0000000000111001};
      array[{4'h1, 4'h3}] = {5'd8, 16'b0000000011110110};
      array[{4'h1, 4'h4}] = {5'd9, 16'b0000000111110101};
      array[{4'h1, 4'h5}] = {5'd11, 16'b0000011111110110};
      array[{4'h1, 4'h6}] = {5'd12, 16'b0000111111110101};
      array[{4'h1, 4'h7}] = {5'd16, 16'b1111111110001000};
      array[{4'h1, 4'h8}] = {5'd16, 16'b1111111110001001};
      array[{4'h1, 4'h9}] = {5'd16, 16'b1111111110001010};
      array[{4'h1, 4'hA}] = {5'd16, 16'b1111111110001011};
      array[{4'h2, 4'h1}] = {5'd5, 16'b0000000000011010};
      array[{4'h2, 4'h2}] = {5'd8, 16'b0000000011110111};
      array[{4'h2, 4'h3}] = {5'd10, 16'b0000001111110111};
      array[{4'h2, 4'h4}] = {5'd12, 16'b0000111111110110};
      array[{4'h2, 4'h5}] = {5'd15, 16'b0111111111000010};
      array[{4'h2, 4'h6}] = {5'd16, 16'b1111111110001100};
      array[{4'h2, 4'h7}] = {5'd16, 16'b1111111110001101};
      array[{4'h2, 4'h8}] = {5'd16, 16'b1111111110001110};
      array[{4'h2, 4'h9}] = {5'd16, 16'b1111111110001111};
      array[{4'h2, 4'hA}] = {5'd16, 16'b1111111110010000};
      array[{4'h3, 4'h1}] = {5'd5, 16'b0000000000011011};
      array[{4'h3, 4'h2}] = {5'd8, 16'b0000000011111000};
      array[{4'h3, 4'h3}] = {5'd10, 16'b0000001111111000};
      array[{4'h3, 4'h4}] = {5'd12, 16'b0000111111110111};
      array[{4'h3, 4'h5}] = {5'd16, 16'b1111111110010001};
      array[{4'h3, 4'h6}] = {5'd16, 16'b1111111110010010};
      array[{4'h3, 4'h7}] = {5'd16, 16'b1111111110010011};
      array[{4'h3, 4'h8}] = {5'd16, 16'b1111111110010100};
      array[{4'h3, 4'h9}] = {5'd16, 16'b1111111110010101};
      array[{4'h3, 4'hA}] = {5'd16, 16'b1111111110010110};
      array[{4'h4, 4'h1}] = {5'd6, 16'b0000000000111010};
      array[{4'h4, 4'h2}] = {5'd9, 16'b0000000111110110};
      array[{4'h4, 4'h3}] = {5'd16, 16'b1111111110010111};
      array[{4'h4, 4'h4}] = {5'd16, 16'b1111111110011000};
      array[{4'h4, 4'h5}] = {5'd16, 16'b1111111110011001};
      array[{4'h4, 4'h6}] = {5'd16, 16'b1111111110011010};
      array[{4'h4, 4'h7}] = {5'd16, 16'b1111111110011011};
      array[{4'h4, 4'h8}] = {5'd16, 16'b1111111110011100};
      array[{4'h4, 4'h9}] = {5'd16, 16'b1111111110011101};
      array[{4'h4, 4'hA}] = {5'd16, 16'b1111111110011110};
      array[{4'h5, 4'h1}] = {5'd6, 16'b0000000000111011};
      array[{4'h5, 4'h2}] = {5'd10, 16'b0000001111111001};
      array[{4'h5, 4'h3}] = {5'd16, 16'b1111111110011111};
      array[{4'h5, 4'h4}] = {5'd16, 16'b1111111110100000};
      array[{4'h5, 4'h5}] = {5'd16, 16'b1111111110100001};
      array[{4'h5, 4'h6}] = {5'd16, 16'b1111111110100010};
      array[{4'h5, 4'h7}] = {5'd16, 16'b1111111110100011};
      array[{4'h5, 4'h8}] = {5'd16, 16'b1111111110100100};
      array[{4'h5, 4'h9}] = {5'd16, 16'b1111111110100101};
      array[{4'h5, 4'hA}] = {5'd16, 16'b1111111110100110};
      array[{4'h6, 4'h1}] = {5'd7, 16'b0000000001111001};
      array[{4'h6, 4'h2}] = {5'd11, 16'b0000011111110111};
      array[{4'h6, 4'h3}] = {5'd16, 16'b1111111110100111};
      array[{4'h6, 4'h4}] = {5'd16, 16'b1111111110101000};
      array[{4'h6, 4'h5}] = {5'd16, 16'b1111111110101001};
      array[{4'h6, 4'h6}] = {5'd16, 16'b1111111110101010};
      array[{4'h6, 4'h7}] = {5'd16, 16'b1111111110101011};
      array[{4'h6, 4'h8}] = {5'd16, 16'b1111111110101100};
      array[{4'h6, 4'h9}] = {5'd16, 16'b1111111110101101};
      array[{4'h6, 4'hA}] = {5'd16, 16'b1111111110101110};
      array[{4'h7, 4'h1}] = {5'd7, 16'b0000000001111010};
      array[{4'h7, 4'h2}] = {5'd11, 16'b0000011111111000};
      array[{4'h7, 4'h3}] = {5'd16, 16'b1111111110101111};
      array[{4'h7, 4'h4}] = {5'd16, 16'b1111111110110000};
      array[{4'h7, 4'h5}] = {5'd16, 16'b1111111110110001};
      array[{4'h7, 4'h6}] = {5'd16, 16'b1111111110110010};
      array[{4'h7, 4'h7}] = {5'd16, 16'b1111111110110011};
      array[{4'h7, 4'h8}] = {5'd16, 16'b1111111110110100};
      array[{4'h7, 4'h9}] = {5'd16, 16'b1111111110110101};
      array[{4'h7, 4'hA}] = {5'd16, 16'b1111111110110110};
      array[{4'h8, 4'h1}] = {5'd8, 16'b0000000011111001};
      array[{4'h8, 4'h2}] = {5'd16, 16'b1111111110110111};
      array[{4'h8, 4'h3}] = {5'd16, 16'b1111111110111000};
      array[{4'h8, 4'h4}] = {5'd16, 16'b1111111110111001};
      array[{4'h8, 4'h5}] = {5'd16, 16'b1111111110111010};
      array[{4'h8, 4'h6}] = {5'd16, 16'b1111111110111011};
      array[{4'h8, 4'h7}] = {5'd16, 16'b1111111110111100};
      array[{4'h8, 4'h8}] = {5'd16, 16'b1111111110111101};
      array[{4'h8, 4'h9}] = {5'd16, 16'b1111111110111110};
      array[{4'h8, 4'hA}] = {5'd16, 16'b1111111110111111};
      array[{4'h9, 4'h1}] = {5'd9, 16'b0000000111110111};
      array[{4'h9, 4'h2}] = {5'd16, 16'b1111111111000000};
      array[{4'h9, 4'h3}] = {5'd16, 16'b1111111111000001};
      array[{4'h9, 4'h4}] = {5'd16, 16'b1111111111000010};
      array[{4'h9, 4'h5}] = {5'd16, 16'b1111111111000011};
      array[{4'h9, 4'h6}] = {5'd16, 16'b1111111111000100};
      array[{4'h9, 4'h7}] = {5'd16, 16'b1111111111000101};
      array[{4'h9, 4'h8}] = {5'd16, 16'b1111111111000110};
      array[{4'h9, 4'h9}] = {5'd16, 16'b1111111111000111};
      array[{4'h9, 4'hA}] = {5'd16, 16'b1111111111001000};
      array[{4'hA, 4'h1}] = {5'd9, 16'b0000000111111000};
      array[{4'hA, 4'h2}] = {5'd16, 16'b1111111111001001};
      array[{4'hA, 4'h3}] = {5'd16, 16'b1111111111001010};
      array[{4'hA, 4'h4}] = {5'd16, 16'b1111111111001011};
      array[{4'hA, 4'h5}] = {5'd16, 16'b1111111111001100};
      array[{4'hA, 4'h6}] = {5'd16, 16'b1111111111001101};
      array[{4'hA, 4'h7}] = {5'd16, 16'b1111111111001110};
      array[{4'hA, 4'h8}] = {5'd16, 16'b1111111111001111};
      array[{4'hA, 4'h9}] = {5'd16, 16'b1111111111010000};
      array[{4'hA, 4'hA}] = {5'd16, 16'b1111111111010001};
      array[{4'hB, 4'h1}] = {5'd9, 16'b0000000111111001};
      array[{4'hB, 4'h2}] = {5'd16, 16'b1111111111010010};
      array[{4'hB, 4'h3}] = {5'd16, 16'b1111111111010011};
      array[{4'hB, 4'h4}] = {5'd16, 16'b1111111111010100};
      array[{4'hB, 4'h5}] = {5'd16, 16'b1111111111010101};
      array[{4'hB, 4'h6}] = {5'd16, 16'b1111111111010110};
      array[{4'hB, 4'h7}] = {5'd16, 16'b1111111111010111};
      array[{4'hB, 4'h8}] = {5'd16, 16'b1111111111011000};
      array[{4'hB, 4'h9}] = {5'd16, 16'b1111111111011001};
      array[{4'hB, 4'hA}] = {5'd16, 16'b1111111111011010};
      array[{4'hC, 4'h1}] = {5'd9, 16'b0000000111111010};
      array[{4'hC, 4'h2}] = {5'd16, 16'b1111111111011011};
      array[{4'hC, 4'h3}] = {5'd16, 16'b1111111111011100};
      array[{4'hC, 4'h4}] = {5'd16, 16'b1111111111011101};
      array[{4'hC, 4'h5}] = {5'd16, 16'b1111111111011110};
      array[{4'hC, 4'h6}] = {5'd16, 16'b1111111111011111};
      array[{4'hC, 4'h7}] = {5'd16, 16'b1111111111100000};
      array[{4'hC, 4'h8}] = {5'd16, 16'b1111111111100001};
      array[{4'hC, 4'h9}] = {5'd16, 16'b1111111111100010};
      array[{4'hC, 4'hA}] = {5'd16, 16'b1111111111100011};
      array[{4'hD, 4'h1}] = {5'd11, 16'b0000011111111001};
      array[{4'hD, 4'h2}] = {5'd16, 16'b1111111111100100};
      array[{4'hD, 4'h3}] = {5'd16, 16'b1111111111100101};
      array[{4'hD, 4'h4}] = {5'd16, 16'b1111111111100110};
      array[{4'hD, 4'h5}] = {5'd16, 16'b1111111111100111};
      array[{4'hD, 4'h6}] = {5'd16, 16'b1111111111101000};
      array[{4'hD, 4'h7}] = {5'd16, 16'b1111111111101001};
      array[{4'hD, 4'h8}] = {5'd16, 16'b1111111111101010};
      array[{4'hD, 4'h9}] = {5'd16, 16'b1111111111101011};
      array[{4'hD, 4'hA}] = {5'd16, 16'b1111111111101100};
      array[{4'hE, 4'h1}] = {5'd14, 16'b0011111111100000};
      array[{4'hE, 4'h2}] = {5'd16, 16'b1111111111101101};
      array[{4'hE, 4'h3}] = {5'd16, 16'b1111111111101110};
      array[{4'hE, 4'h4}] = {5'd16, 16'b1111111111101111};
      array[{4'hE, 4'h5}] = {5'd16, 16'b1111111111110000};
      array[{4'hE, 4'h6}] = {5'd16, 16'b1111111111110001};
      array[{4'hE, 4'h7}] = {5'd16, 16'b1111111111110010};
      array[{4'hE, 4'h8}] = {5'd16, 16'b1111111111110011};
      array[{4'hE, 4'h9}] = {5'd16, 16'b1111111111110100};
      array[{4'hE, 4'hA}] = {5'd16, 16'b1111111111110101};
      array[{4'hF, 4'h0}] = {5'd10, 16'b0000001111111010};
      array[{4'hF, 4'h1}] = {5'd15, 16'b0111111111000011};
      array[{4'hF, 4'h2}] = {5'd16, 16'b1111111111110110};
      array[{4'hF, 4'h3}] = {5'd16, 16'b1111111111110111};
      array[{4'hF, 4'h4}] = {5'd16, 16'b1111111111111000};
      array[{4'hF, 4'h5}] = {5'd16, 16'b1111111111111001};
      array[{4'hF, 4'h6}] = {5'd16, 16'b1111111111111010};
      array[{4'hF, 4'h7}] = {5'd16, 16'b1111111111111011};
      array[{4'hF, 4'h8}] = {5'd16, 16'b1111111111111100};
      array[{4'hF, 4'h9}] = {5'd16, 16'b1111111111111101};
      array[{4'hF, 4'hA}] = {5'd16, 16'b1111111111111110};
    end
end
endmodule
